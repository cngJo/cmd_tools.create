module main

fn main() {
    println('create')
}